module reg32(); 
endmodule